`timescale 1 ps / 1 ps
module letter(
	input [7:0] number,
	output reg [19:0] digit [0:5]
);

	always @* begin
		case (number)
			7'd71: begin // G
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000000000;
				digit[3] = 20'b11111000001111111111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			7'd69: begin // E
				digit[0] = 20'b11111111111111111111;
				digit[1] = 20'b11111000000000000000;
				digit[2] = 20'b11111111111111100000;
				digit[3] = 20'b11111000000000000000;
				digit[4] = 20'b11111000000000000000;
				digit[5] = 20'b11111111111111111111;
			end
			
			7'd83: begin // S
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b00000111110000000000;
				digit[3] = 20'b00000000001111100000;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			7'd84: begin // T
				digit[0] = 20'b11111111111111111111;
				digit[1] = 20'b00000000001111100000;
				digit[2] = 20'b00000000001111100000;
				digit[3] = 20'b00000000001111100000;
				digit[4] = 20'b00000000001111100000;
				digit[5] = 20'b00000000001111100000;
			end
			
			7'd85: begin // U
				digit[0] = 20'b11111000000000011111;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			7'd82: begin // R
				digit[0] = 20'b11111111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111111111111100000;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b11111000000000011111;
			end
			
			7'd65: begin // A
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111111111111111111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b11111000000000011111;
			end
			
			7'd80: begin // P
				digit[0] = 20'b11111111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111111111111100000;
				digit[4] = 20'b11111000000000000000;
				digit[5] = 20'b11111000000000000000;
			end
			
			7'd68: begin // D
				digit[0] = 20'b11111111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b11111111111111100000;
			end
		endcase
	end

endmodule