`timescale 1 ps / 1 ps
module digit(
	input [3:0] number,
	output reg [19:0] digit [0:5]
);

	always @* begin
		case (number)
			4'd0: begin
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			4'd1: begin
				digit[0] = 20'b00000000001111100000;
				digit[1] = 20'b00000111111111100000;
				digit[2] = 20'b11111000001111100000;
				digit[3] = 20'b00000000001111100000;
				digit[4] = 20'b00000000001111100000;
				digit[5] = 20'b11111111111111111111;
			end
			
			4'd2: begin
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b00000000000000011111;
				digit[3] = 20'b00000111111111100000;
				digit[4] = 20'b11111000000000000000;
				digit[5] = 20'b11111111111111111111;
			end
			
			4'd3: begin
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b00000000001111100000;
				digit[3] = 20'b00000000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			4'd4: begin
				digit[0] = 20'b00000000001111111111;
				digit[1] = 20'b00000111110000011111;
				digit[2] = 20'b11111000000000011111;
				digit[3] = 20'b11111111111111111111;
				digit[4] = 20'b00000000000000011111;
				digit[5] = 20'b00000000000000011111;
			end
			
			4'd5: begin
				digit[0] = 20'b11111111111111111111;
				digit[1] = 20'b11111000000000000000;
				digit[2] = 20'b11111111111111100000;
				digit[3] = 20'b00000000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			4'd6: begin
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b11111000000000000000;
				digit[3] = 20'b11111111111111100000;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			4'd7: begin
				digit[0] = 20'b11111111111111111111;
				digit[1] = 20'b00000000000000011111;
				digit[2] = 20'b00000000001111100000;
				digit[3] = 20'b00000111110000000000;
				digit[4] = 20'b11111000000000000000;
				digit[5] = 20'b11111000000000000000;
			end
			
			4'd8: begin
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b00000111111111100000;
				digit[3] = 20'b11111000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end
			
			4'd9: begin
				digit[0] = 20'b00000111111111100000;
				digit[1] = 20'b11111000000000011111;
				digit[2] = 20'b00000111111111111111;
				digit[3] = 20'b00000000000000011111;
				digit[4] = 20'b11111000000000011111;
				digit[5] = 20'b00000111111111100000;
			end

		endcase
	end

endmodule