`timescale 1 ps / 1 ps
module digit(
	input [3:0] number,
	output reg [29:0] digit [0:3]
);

	always @* begin
		case (number)
			4'd0: begin
				digit[0] = 30'b000001111111111111111111100000;
				digit[1] = 30'b111110000000000000000000011111;
				digit[2] = 30'b111110000000000000000000011111;
				digit[3] = 30'b000001111111111111111111100000;
			end
			
			4'd1: begin
				digit[0] = 30'b111110000000000111110000000000;
				digit[1] = 30'b111110000000000000001111100000;
				digit[2] = 30'b111111111111111111111111111111;
				digit[3] = 30'b111110000000000000000000000000;
			end
				
			4'd2: begin
				digit[0] = 30'b111111111100000000001111100000;
				digit[1] = 30'b111110000011111000000000011111;
				digit[2] = 30'b111110000011111000000000011111;
				digit[3] = 30'b111110000000000111111111100000;
			end
				
			4'd3: begin
				digit[0] = 30'b000001111100000000001111100000;
				digit[1] = 30'b111110000000000000000000011111;
				digit[2] = 30'b111110000000000111110000011111;
				digit[3] = 30'b000001111111111000001111100000;
			end
			
			4'd4: begin
				digit[0] = 30'b000000000011111111110000000000;
				digit[1] = 30'b000000000011111000001111100000;
				digit[2] = 30'b000000000011111000000000011111;
				digit[3] = 30'b111111111111111111111111111111;
			end
			
			4'd5: begin
				digit[0] = 30'b000001111100000111111111111111;
				digit[1] = 30'b111110000000000111110000011111;
				digit[2] = 30'b111110000000000111110000011111;
				digit[3] = 30'b000001111111111000000000011111;
			end
				
			4'd6: begin
				digit[0] = 30'b000001111111111111111111100000;
				digit[1] = 30'b111110000011111000000000011111;
				digit[2] = 30'b111110000011111000000000011111;
				digit[3] = 30'b000001111100000000001111100000;
			end
				
			4'd7: begin
				digit[0] = 30'b111111111100000000000000011111;
				digit[1] = 30'b000000000011111000000000011111;
				digit[2] = 30'b000000000000000111110000011111;
				digit[3] = 30'b000000000000000000001111111111;
			end
				
			4'd8: begin
				digit[0] = 30'b000001111111111000001111100000;
				digit[1] = 30'b111110000000000111110000011111;
				digit[2] = 30'b111110000000000111110000011111;
				digit[3] = 30'b000001111111111000001111100000;
			end
				
			4'd9: begin
				digit[0] = 30'b000001111100000000001111100000;
				digit[1] = 30'b111110000000000111110000011111;
				digit[2] = 30'b111110000000000111110000011111;
				digit[3] = 30'b000001111111111111111111100000;
			end
				

		endcase
	end

endmodule