`timescale 1 ps / 1 ps
module letter(
	input [7:0] number,
	output reg [29:0] digit [0:3]
);

	always @* begin
		case (number)
			7'd88: begin // X
				digit[0] = 30'b000000000000000000000000000000;
				digit[1] = 30'b111111111111111000001111111111;
				digit[2] = 30'b000000000000000111110000000000;
				digit[3] = 30'b111111111111111000001111111111;
			end
			
			7'd89: begin // Y
				digit[0] = 30'b000000000000000000000000000000;
				digit[1] = 30'b000000000000000111111111111111;
				digit[2] = 30'b111111111111111000000000000000;
				digit[3] = 30'b000000000000000111111111111111;
			end
			
			7'd84: begin // T
				digit[0] = 30'b000000000000000000000000000000;
				digit[1] = 30'b000000000000000000000000011111;
				digit[2] = 30'b111111111111111111111111111111;
				digit[3] = 30'b000000000000000000000000011111;
			end
			
			7'd65: begin // A
				digit[0] = 30'b111111111111111111111111100000;
				digit[1] = 30'b000000000011111000000000011111;
				digit[2] = 30'b000000000011111000000000011111;
				digit[3] = 30'b111111111111111111111111100000;
			end
			
			7'd80: begin // P
				digit[0] = 30'b111111111111111111111111111111;
				digit[1] = 30'b000000000011111000000000011111;
				digit[2] = 30'b000000000011111000000000011111;
				digit[3] = 30'b000000000000000111111111100000;
			end
			
			7'd68: begin // D
				digit[0] = 30'b111111111111111111111111111111;
				digit[1] = 30'b111110000000000000000000011111;
				digit[2] = 30'b111110000000000000000000011111;
				digit[3] = 30'b000001111111111111111111100000;
			end
			
			7'd82: begin // R
				digit[0] = 30'b111111111111111111111111111111;
				digit[1] = 30'b000000000011111000000000011111;
				digit[2] = 30'b000000000011111000000000011111;
				digit[3] = 30'b111111111100000111111111100000;
			end
			
			7'd71: begin // G
				digit[0] = 30'b000001111111111111111111100000;
				digit[1] = 30'b111110000000000000000000011111;
				digit[2] = 30'b111110000011111000000000011111;
				digit[3] = 30'b000001111111111000001111100000;
			end
			
			7'd73: begin // I
				digit[0] = 30'b000000000000000000000000000000;
				digit[1] = 30'b111110000000000000000000011111;
				digit[2] = 30'b111111111111111111111111111111;
				digit[3] = 30'b111110000000000000000000011111;
			end
			
			7'd76: begin // L
				digit[0] = 30'b111111111111111111111111111111;
				digit[1] = 30'b111110000000000000000000000000;
				digit[2] = 30'b111110000000000000000000000000;
				digit[3] = 30'b111110000000000000000000000000;
			end
			
			7'd69: begin // E
				digit[0] = 30'b111111111111111111111111111111;
				digit[1] = 30'b111110000000000111110000011111;
				digit[2] = 30'b111110000000000111110000011111;
				digit[3] = 30'b111110000000000000000000011111;
			end
			
		endcase
	end

endmodule